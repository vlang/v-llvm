module vllvm

import bindings

pub const (
	version = '0.1.0'
)